LINJARA KOMPONENTER, RESISTANS - UPPGIFT 1.4.1

.OPTIONS POST

R1 IN 0 3.3K
IIN 0 IN 1M

.DC IIN 0 1M 0.1M

.END

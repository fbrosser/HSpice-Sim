ICKELINJARA KOMPONENTER, DIOD - UPPGIFT 1.4.2

.OPTIONS POST

.MODEL DIOD D LEVEL=1 IS=1F

D1 IN 0 DIOD
IIN 0 IN 1M

.DC IIN 0 1M 0.01M

.END

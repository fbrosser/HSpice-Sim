J-OMEGA-Metoden - UPPGIFT 1.5.1

.OPTIONS POST

.MODEL DIOD D LEVEL=1 IS=1F

R1 IN UT 3.3K
C1 UT 0 1N
VIN IN 0 SIN(0 1 10K)

.TRAN 0.01U 1M

.END

I-V SIMULERING AV LASTRESISTANS

.PARAM SUPPLYV=3.3V
.OPTIONS POST

R2 VDD UT 15000

VVDD VDD 0 DC SUPPLYV
VUT UT 0 DC SUPPLYV

.DC VUT 0 SUPPLYV 0.1

.PROBE IR2=PAR('-I(VVDD)')

.END

SIMULERING AV SPANNINGSDELNING OVER RESISTANSER - UPPGIFT 1.3.3

.PARAM SUPPLYV=3.3

.OPTIONS POST

R1 VDD UT 3300
R2 UT 0 10K

VVDD VDD 0 DC SUPPLYV

.TRAN 0.1U 1M

.END
